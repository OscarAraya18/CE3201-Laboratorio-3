module CompuertaOR(operandoA, operandoB, resultado);
	parameter ancho = 'd3;
	input [ancho:0] operandoA;
	input [ancho:0] operandoB;
	output [ancho:0] resultado;
	assign resultado = operandoA | operandoB;
endmodule 