module DetectorCero #(parameter ancho = 'd3) (operandoA, operandoB, resultado, carryOut);


endmodule 